// Sigmoid Function using a LUT
`timescale 1ns / 1ps


module sigmoid
#(
    parameter Q = 13,   // Fractional part
    parameter N = 16, 
    parameter MEM_SIZE = 10 
)
(
    input          clk,
    input          rstn,
    input    [N-1:0] sigmoid_in,
    output   [N-1:0] sigmoid_out
);

// Note: To save space, we are truncating extra decimal points 

// Load the memory file
reg [N-1:0] sigmoid_mem [0:2**MEM_SIZE-1];
wire [MEM_SIZE-1:0] x_trunc; 
assign x_trunc = sigmoid_in[N-1:N-MEM_SIZE];
reg [MEM_SIZE-1:0] y;

// ----------- AUTOGENERATED CODE -------------------------- // 
assign sigmoid_mem[0] = 16'b0000000010010100;
assign sigmoid_mem[1] = 16'b0000000010010101;
assign sigmoid_mem[2] = 16'b0000000010010110;
assign sigmoid_mem[3] = 16'b0000000010010111;
assign sigmoid_mem[4] = 16'b0000000010011001;
assign sigmoid_mem[5] = 16'b0000000010011010;
assign sigmoid_mem[6] = 16'b0000000010011011;
assign sigmoid_mem[7] = 16'b0000000010011100;
assign sigmoid_mem[8] = 16'b0000000010011101;
assign sigmoid_mem[9] = 16'b0000000010011111;
assign sigmoid_mem[10] = 16'b0000000010100000;
assign sigmoid_mem[11] = 16'b0000000010100001;
assign sigmoid_mem[12] = 16'b0000000010100010;
assign sigmoid_mem[13] = 16'b0000000010100100;
assign sigmoid_mem[14] = 16'b0000000010100101;
assign sigmoid_mem[15] = 16'b0000000010100110;
assign sigmoid_mem[16] = 16'b0000000010100111;
assign sigmoid_mem[17] = 16'b0000000010101001;
assign sigmoid_mem[18] = 16'b0000000010101010;
assign sigmoid_mem[19] = 16'b0000000010101011;
assign sigmoid_mem[20] = 16'b0000000010101101;
assign sigmoid_mem[21] = 16'b0000000010101110;
assign sigmoid_mem[22] = 16'b0000000010101111;
assign sigmoid_mem[23] = 16'b0000000010110001;
assign sigmoid_mem[24] = 16'b0000000010110010;
assign sigmoid_mem[25] = 16'b0000000010110011;
assign sigmoid_mem[26] = 16'b0000000010110101;
assign sigmoid_mem[27] = 16'b0000000010110110;
assign sigmoid_mem[28] = 16'b0000000010110111;
assign sigmoid_mem[29] = 16'b0000000010111001;
assign sigmoid_mem[30] = 16'b0000000010111010;
assign sigmoid_mem[31] = 16'b0000000010111100;
assign sigmoid_mem[32] = 16'b0000000010111101;
assign sigmoid_mem[33] = 16'b0000000010111111;
assign sigmoid_mem[34] = 16'b0000000011000000;
assign sigmoid_mem[35] = 16'b0000000011000010;
assign sigmoid_mem[36] = 16'b0000000011000011;
assign sigmoid_mem[37] = 16'b0000000011000101;
assign sigmoid_mem[38] = 16'b0000000011000110;
assign sigmoid_mem[39] = 16'b0000000011001000;
assign sigmoid_mem[40] = 16'b0000000011001001;
assign sigmoid_mem[41] = 16'b0000000011001011;
assign sigmoid_mem[42] = 16'b0000000011001100;
assign sigmoid_mem[43] = 16'b0000000011001110;
assign sigmoid_mem[44] = 16'b0000000011001111;
assign sigmoid_mem[45] = 16'b0000000011010001;
assign sigmoid_mem[46] = 16'b0000000011010011;
assign sigmoid_mem[47] = 16'b0000000011010100;
assign sigmoid_mem[48] = 16'b0000000011010110;
assign sigmoid_mem[49] = 16'b0000000011010111;
assign sigmoid_mem[50] = 16'b0000000011011001;
assign sigmoid_mem[51] = 16'b0000000011011011;
assign sigmoid_mem[52] = 16'b0000000011011100;
assign sigmoid_mem[53] = 16'b0000000011011110;
assign sigmoid_mem[54] = 16'b0000000011100000;
assign sigmoid_mem[55] = 16'b0000000011100001;
assign sigmoid_mem[56] = 16'b0000000011100011;
assign sigmoid_mem[57] = 16'b0000000011100101;
assign sigmoid_mem[58] = 16'b0000000011100111;
assign sigmoid_mem[59] = 16'b0000000011101000;
assign sigmoid_mem[60] = 16'b0000000011101010;
assign sigmoid_mem[61] = 16'b0000000011101100;
assign sigmoid_mem[62] = 16'b0000000011101110;
assign sigmoid_mem[63] = 16'b0000000011110000;
assign sigmoid_mem[64] = 16'b0000000011110001;
assign sigmoid_mem[65] = 16'b0000000011110011;
assign sigmoid_mem[66] = 16'b0000000011110101;
assign sigmoid_mem[67] = 16'b0000000011110111;
assign sigmoid_mem[68] = 16'b0000000011111001;
assign sigmoid_mem[69] = 16'b0000000011111011;
assign sigmoid_mem[70] = 16'b0000000011111101;
assign sigmoid_mem[71] = 16'b0000000011111111;
assign sigmoid_mem[72] = 16'b0000000100000001;
assign sigmoid_mem[73] = 16'b0000000100000011;
assign sigmoid_mem[74] = 16'b0000000100000100;
assign sigmoid_mem[75] = 16'b0000000100000110;
assign sigmoid_mem[76] = 16'b0000000100001000;
assign sigmoid_mem[77] = 16'b0000000100001010;
assign sigmoid_mem[78] = 16'b0000000100001101;
assign sigmoid_mem[79] = 16'b0000000100001111;
assign sigmoid_mem[80] = 16'b0000000100010001;
assign sigmoid_mem[81] = 16'b0000000100010011;
assign sigmoid_mem[82] = 16'b0000000100010101;
assign sigmoid_mem[83] = 16'b0000000100010111;
assign sigmoid_mem[84] = 16'b0000000100011001;
assign sigmoid_mem[85] = 16'b0000000100011011;
assign sigmoid_mem[86] = 16'b0000000100011101;
assign sigmoid_mem[87] = 16'b0000000100011111;
assign sigmoid_mem[88] = 16'b0000000100100010;
assign sigmoid_mem[89] = 16'b0000000100100100;
assign sigmoid_mem[90] = 16'b0000000100100110;
assign sigmoid_mem[91] = 16'b0000000100101000;
assign sigmoid_mem[92] = 16'b0000000100101010;
assign sigmoid_mem[93] = 16'b0000000100101101;
assign sigmoid_mem[94] = 16'b0000000100101111;
assign sigmoid_mem[95] = 16'b0000000100110001;
assign sigmoid_mem[96] = 16'b0000000100110100;
assign sigmoid_mem[97] = 16'b0000000100110110;
assign sigmoid_mem[98] = 16'b0000000100111000;
assign sigmoid_mem[99] = 16'b0000000100111011;
assign sigmoid_mem[100] = 16'b0000000100111101;
assign sigmoid_mem[101] = 16'b0000000100111111;
assign sigmoid_mem[102] = 16'b0000000101000010;
assign sigmoid_mem[103] = 16'b0000000101000100;
assign sigmoid_mem[104] = 16'b0000000101000111;
assign sigmoid_mem[105] = 16'b0000000101001001;
assign sigmoid_mem[106] = 16'b0000000101001100;
assign sigmoid_mem[107] = 16'b0000000101001110;
assign sigmoid_mem[108] = 16'b0000000101010001;
assign sigmoid_mem[109] = 16'b0000000101010011;
assign sigmoid_mem[110] = 16'b0000000101010110;
assign sigmoid_mem[111] = 16'b0000000101011000;
assign sigmoid_mem[112] = 16'b0000000101011011;
assign sigmoid_mem[113] = 16'b0000000101011101;
assign sigmoid_mem[114] = 16'b0000000101100000;
assign sigmoid_mem[115] = 16'b0000000101100011;
assign sigmoid_mem[116] = 16'b0000000101100101;
assign sigmoid_mem[117] = 16'b0000000101101000;
assign sigmoid_mem[118] = 16'b0000000101101011;
assign sigmoid_mem[119] = 16'b0000000101101110;
assign sigmoid_mem[120] = 16'b0000000101110000;
assign sigmoid_mem[121] = 16'b0000000101110011;
assign sigmoid_mem[122] = 16'b0000000101110110;
assign sigmoid_mem[123] = 16'b0000000101111001;
assign sigmoid_mem[124] = 16'b0000000101111011;
assign sigmoid_mem[125] = 16'b0000000101111110;
assign sigmoid_mem[126] = 16'b0000000110000001;
assign sigmoid_mem[127] = 16'b0000000110000100;
assign sigmoid_mem[128] = 16'b0000000110000111;
assign sigmoid_mem[129] = 16'b0000000110001010;
assign sigmoid_mem[130] = 16'b0000000110001101;
assign sigmoid_mem[131] = 16'b0000000110010000;
assign sigmoid_mem[132] = 16'b0000000110010011;
assign sigmoid_mem[133] = 16'b0000000110010110;
assign sigmoid_mem[134] = 16'b0000000110011001;
assign sigmoid_mem[135] = 16'b0000000110011100;
assign sigmoid_mem[136] = 16'b0000000110011111;
assign sigmoid_mem[137] = 16'b0000000110100010;
assign sigmoid_mem[138] = 16'b0000000110100101;
assign sigmoid_mem[139] = 16'b0000000110101000;
assign sigmoid_mem[140] = 16'b0000000110101011;
assign sigmoid_mem[141] = 16'b0000000110101111;
assign sigmoid_mem[142] = 16'b0000000110110010;
assign sigmoid_mem[143] = 16'b0000000110110101;
assign sigmoid_mem[144] = 16'b0000000110111000;
assign sigmoid_mem[145] = 16'b0000000110111011;
assign sigmoid_mem[146] = 16'b0000000110111111;
assign sigmoid_mem[147] = 16'b0000000111000010;
assign sigmoid_mem[148] = 16'b0000000111000101;
assign sigmoid_mem[149] = 16'b0000000111001001;
assign sigmoid_mem[150] = 16'b0000000111001100;
assign sigmoid_mem[151] = 16'b0000000111010000;
assign sigmoid_mem[152] = 16'b0000000111010011;
assign sigmoid_mem[153] = 16'b0000000111010110;
assign sigmoid_mem[154] = 16'b0000000111011010;
assign sigmoid_mem[155] = 16'b0000000111011101;
assign sigmoid_mem[156] = 16'b0000000111100001;
assign sigmoid_mem[157] = 16'b0000000111100101;
assign sigmoid_mem[158] = 16'b0000000111101000;
assign sigmoid_mem[159] = 16'b0000000111101100;
assign sigmoid_mem[160] = 16'b0000000111101111;
assign sigmoid_mem[161] = 16'b0000000111110011;
assign sigmoid_mem[162] = 16'b0000000111110111;
assign sigmoid_mem[163] = 16'b0000000111111010;
assign sigmoid_mem[164] = 16'b0000000111111110;
assign sigmoid_mem[165] = 16'b0000001000000010;
assign sigmoid_mem[166] = 16'b0000001000000110;
assign sigmoid_mem[167] = 16'b0000001000001001;
assign sigmoid_mem[168] = 16'b0000001000001101;
assign sigmoid_mem[169] = 16'b0000001000010001;
assign sigmoid_mem[170] = 16'b0000001000010101;
assign sigmoid_mem[171] = 16'b0000001000011001;
assign sigmoid_mem[172] = 16'b0000001000011101;
assign sigmoid_mem[173] = 16'b0000001000100001;
assign sigmoid_mem[174] = 16'b0000001000100101;
assign sigmoid_mem[175] = 16'b0000001000101001;
assign sigmoid_mem[176] = 16'b0000001000101101;
assign sigmoid_mem[177] = 16'b0000001000110001;
assign sigmoid_mem[178] = 16'b0000001000110101;
assign sigmoid_mem[179] = 16'b0000001000111001;
assign sigmoid_mem[180] = 16'b0000001000111101;
assign sigmoid_mem[181] = 16'b0000001001000010;
assign sigmoid_mem[182] = 16'b0000001001000110;
assign sigmoid_mem[183] = 16'b0000001001001010;
assign sigmoid_mem[184] = 16'b0000001001001110;
assign sigmoid_mem[185] = 16'b0000001001010011;
assign sigmoid_mem[186] = 16'b0000001001010111;
assign sigmoid_mem[187] = 16'b0000001001011011;
assign sigmoid_mem[188] = 16'b0000001001100000;
assign sigmoid_mem[189] = 16'b0000001001100100;
assign sigmoid_mem[190] = 16'b0000001001101000;
assign sigmoid_mem[191] = 16'b0000001001101101;
assign sigmoid_mem[192] = 16'b0000001001110001;
assign sigmoid_mem[193] = 16'b0000001001110110;
assign sigmoid_mem[194] = 16'b0000001001111011;
assign sigmoid_mem[195] = 16'b0000001001111111;
assign sigmoid_mem[196] = 16'b0000001010000100;
assign sigmoid_mem[197] = 16'b0000001010001000;
assign sigmoid_mem[198] = 16'b0000001010001101;
assign sigmoid_mem[199] = 16'b0000001010010010;
assign sigmoid_mem[200] = 16'b0000001010010111;
assign sigmoid_mem[201] = 16'b0000001010011011;
assign sigmoid_mem[202] = 16'b0000001010100000;
assign sigmoid_mem[203] = 16'b0000001010100101;
assign sigmoid_mem[204] = 16'b0000001010101010;
assign sigmoid_mem[205] = 16'b0000001010101111;
assign sigmoid_mem[206] = 16'b0000001010110100;
assign sigmoid_mem[207] = 16'b0000001010111001;
assign sigmoid_mem[208] = 16'b0000001010111110;
assign sigmoid_mem[209] = 16'b0000001011000011;
assign sigmoid_mem[210] = 16'b0000001011001000;
assign sigmoid_mem[211] = 16'b0000001011001101;
assign sigmoid_mem[212] = 16'b0000001011010010;
assign sigmoid_mem[213] = 16'b0000001011010111;
assign sigmoid_mem[214] = 16'b0000001011011100;
assign sigmoid_mem[215] = 16'b0000001011100010;
assign sigmoid_mem[216] = 16'b0000001011100111;
assign sigmoid_mem[217] = 16'b0000001011101100;
assign sigmoid_mem[218] = 16'b0000001011110001;
assign sigmoid_mem[219] = 16'b0000001011110111;
assign sigmoid_mem[220] = 16'b0000001011111100;
assign sigmoid_mem[221] = 16'b0000001100000010;
assign sigmoid_mem[222] = 16'b0000001100000111;
assign sigmoid_mem[223] = 16'b0000001100001101;
assign sigmoid_mem[224] = 16'b0000001100010010;
assign sigmoid_mem[225] = 16'b0000001100011000;
assign sigmoid_mem[226] = 16'b0000001100011101;
assign sigmoid_mem[227] = 16'b0000001100100011;
assign sigmoid_mem[228] = 16'b0000001100101001;
assign sigmoid_mem[229] = 16'b0000001100101110;
assign sigmoid_mem[230] = 16'b0000001100110100;
assign sigmoid_mem[231] = 16'b0000001100111010;
assign sigmoid_mem[232] = 16'b0000001101000000;
assign sigmoid_mem[233] = 16'b0000001101000110;
assign sigmoid_mem[234] = 16'b0000001101001011;
assign sigmoid_mem[235] = 16'b0000001101010001;
assign sigmoid_mem[236] = 16'b0000001101010111;
assign sigmoid_mem[237] = 16'b0000001101011101;
assign sigmoid_mem[238] = 16'b0000001101100011;
assign sigmoid_mem[239] = 16'b0000001101101010;
assign sigmoid_mem[240] = 16'b0000001101110000;
assign sigmoid_mem[241] = 16'b0000001101110110;
assign sigmoid_mem[242] = 16'b0000001101111100;
assign sigmoid_mem[243] = 16'b0000001110000010;
assign sigmoid_mem[244] = 16'b0000001110001000;
assign sigmoid_mem[245] = 16'b0000001110001111;
assign sigmoid_mem[246] = 16'b0000001110010101;
assign sigmoid_mem[247] = 16'b0000001110011100;
assign sigmoid_mem[248] = 16'b0000001110100010;
assign sigmoid_mem[249] = 16'b0000001110101000;
assign sigmoid_mem[250] = 16'b0000001110101111;
assign sigmoid_mem[251] = 16'b0000001110110101;
assign sigmoid_mem[252] = 16'b0000001110111100;
assign sigmoid_mem[253] = 16'b0000001111000011;
assign sigmoid_mem[254] = 16'b0000001111001001;
assign sigmoid_mem[255] = 16'b0000001111010000;
assign sigmoid_mem[256] = 16'b0000001111010111;
assign sigmoid_mem[257] = 16'b0000001111011110;
assign sigmoid_mem[258] = 16'b0000001111100100;
assign sigmoid_mem[259] = 16'b0000001111101011;
assign sigmoid_mem[260] = 16'b0000001111110010;
assign sigmoid_mem[261] = 16'b0000001111111001;
assign sigmoid_mem[262] = 16'b0000010000000000;
assign sigmoid_mem[263] = 16'b0000010000000111;
assign sigmoid_mem[264] = 16'b0000010000001110;
assign sigmoid_mem[265] = 16'b0000010000010101;
assign sigmoid_mem[266] = 16'b0000010000011100;
assign sigmoid_mem[267] = 16'b0000010000100100;
assign sigmoid_mem[268] = 16'b0000010000101011;
assign sigmoid_mem[269] = 16'b0000010000110010;
assign sigmoid_mem[270] = 16'b0000010000111001;
assign sigmoid_mem[271] = 16'b0000010001000001;
assign sigmoid_mem[272] = 16'b0000010001001000;
assign sigmoid_mem[273] = 16'b0000010001010000;
assign sigmoid_mem[274] = 16'b0000010001010111;
assign sigmoid_mem[275] = 16'b0000010001011111;
assign sigmoid_mem[276] = 16'b0000010001100110;
assign sigmoid_mem[277] = 16'b0000010001101110;
assign sigmoid_mem[278] = 16'b0000010001110101;
assign sigmoid_mem[279] = 16'b0000010001111101;
assign sigmoid_mem[280] = 16'b0000010010000101;
assign sigmoid_mem[281] = 16'b0000010010001101;
assign sigmoid_mem[282] = 16'b0000010010010100;
assign sigmoid_mem[283] = 16'b0000010010011100;
assign sigmoid_mem[284] = 16'b0000010010100100;
assign sigmoid_mem[285] = 16'b0000010010101100;
assign sigmoid_mem[286] = 16'b0000010010110100;
assign sigmoid_mem[287] = 16'b0000010010111100;
assign sigmoid_mem[288] = 16'b0000010011000100;
assign sigmoid_mem[289] = 16'b0000010011001101;
assign sigmoid_mem[290] = 16'b0000010011010101;
assign sigmoid_mem[291] = 16'b0000010011011101;
assign sigmoid_mem[292] = 16'b0000010011100101;
assign sigmoid_mem[293] = 16'b0000010011101110;
assign sigmoid_mem[294] = 16'b0000010011110110;
assign sigmoid_mem[295] = 16'b0000010011111110;
assign sigmoid_mem[296] = 16'b0000010100000111;
assign sigmoid_mem[297] = 16'b0000010100001111;
assign sigmoid_mem[298] = 16'b0000010100011000;
assign sigmoid_mem[299] = 16'b0000010100100000;
assign sigmoid_mem[300] = 16'b0000010100101001;
assign sigmoid_mem[301] = 16'b0000010100110010;
assign sigmoid_mem[302] = 16'b0000010100111010;
assign sigmoid_mem[303] = 16'b0000010101000011;
assign sigmoid_mem[304] = 16'b0000010101001100;
assign sigmoid_mem[305] = 16'b0000010101010101;
assign sigmoid_mem[306] = 16'b0000010101011110;
assign sigmoid_mem[307] = 16'b0000010101100111;
assign sigmoid_mem[308] = 16'b0000010101110000;
assign sigmoid_mem[309] = 16'b0000010101111001;
assign sigmoid_mem[310] = 16'b0000010110000010;
assign sigmoid_mem[311] = 16'b0000010110001011;
assign sigmoid_mem[312] = 16'b0000010110010100;
assign sigmoid_mem[313] = 16'b0000010110011110;
assign sigmoid_mem[314] = 16'b0000010110100111;
assign sigmoid_mem[315] = 16'b0000010110110000;
assign sigmoid_mem[316] = 16'b0000010110111010;
assign sigmoid_mem[317] = 16'b0000010111000011;
assign sigmoid_mem[318] = 16'b0000010111001100;
assign sigmoid_mem[319] = 16'b0000010111010110;
assign sigmoid_mem[320] = 16'b0000010111011111;
assign sigmoid_mem[321] = 16'b0000010111101001;
assign sigmoid_mem[322] = 16'b0000010111110011;
assign sigmoid_mem[323] = 16'b0000010111111100;
assign sigmoid_mem[324] = 16'b0000011000000110;
assign sigmoid_mem[325] = 16'b0000011000010000;
assign sigmoid_mem[326] = 16'b0000011000011010;
assign sigmoid_mem[327] = 16'b0000011000100100;
assign sigmoid_mem[328] = 16'b0000011000101110;
assign sigmoid_mem[329] = 16'b0000011000111000;
assign sigmoid_mem[330] = 16'b0000011001000010;
assign sigmoid_mem[331] = 16'b0000011001001100;
assign sigmoid_mem[332] = 16'b0000011001010110;
assign sigmoid_mem[333] = 16'b0000011001100000;
assign sigmoid_mem[334] = 16'b0000011001101010;
assign sigmoid_mem[335] = 16'b0000011001110101;
assign sigmoid_mem[336] = 16'b0000011001111111;
assign sigmoid_mem[337] = 16'b0000011010001001;
assign sigmoid_mem[338] = 16'b0000011010010100;
assign sigmoid_mem[339] = 16'b0000011010011110;
assign sigmoid_mem[340] = 16'b0000011010101001;
assign sigmoid_mem[341] = 16'b0000011010110011;
assign sigmoid_mem[342] = 16'b0000011010111110;
assign sigmoid_mem[343] = 16'b0000011011001001;
assign sigmoid_mem[344] = 16'b0000011011010011;
assign sigmoid_mem[345] = 16'b0000011011011110;
assign sigmoid_mem[346] = 16'b0000011011101001;
assign sigmoid_mem[347] = 16'b0000011011110100;
assign sigmoid_mem[348] = 16'b0000011011111111;
assign sigmoid_mem[349] = 16'b0000011100001010;
assign sigmoid_mem[350] = 16'b0000011100010101;
assign sigmoid_mem[351] = 16'b0000011100100000;
assign sigmoid_mem[352] = 16'b0000011100101011;
assign sigmoid_mem[353] = 16'b0000011100110110;
assign sigmoid_mem[354] = 16'b0000011101000001;
assign sigmoid_mem[355] = 16'b0000011101001101;
assign sigmoid_mem[356] = 16'b0000011101011000;
assign sigmoid_mem[357] = 16'b0000011101100011;
assign sigmoid_mem[358] = 16'b0000011101101111;
assign sigmoid_mem[359] = 16'b0000011101111010;
assign sigmoid_mem[360] = 16'b0000011110000110;
assign sigmoid_mem[361] = 16'b0000011110010001;
assign sigmoid_mem[362] = 16'b0000011110011101;
assign sigmoid_mem[363] = 16'b0000011110101000;
assign sigmoid_mem[364] = 16'b0000011110110100;
assign sigmoid_mem[365] = 16'b0000011111000000;
assign sigmoid_mem[366] = 16'b0000011111001011;
assign sigmoid_mem[367] = 16'b0000011111010111;
assign sigmoid_mem[368] = 16'b0000011111100011;
assign sigmoid_mem[369] = 16'b0000011111101111;
assign sigmoid_mem[370] = 16'b0000011111111011;
assign sigmoid_mem[371] = 16'b0000100000000111;
assign sigmoid_mem[372] = 16'b0000100000010011;
assign sigmoid_mem[373] = 16'b0000100000011111;
assign sigmoid_mem[374] = 16'b0000100000101011;
assign sigmoid_mem[375] = 16'b0000100000110111;
assign sigmoid_mem[376] = 16'b0000100001000100;
assign sigmoid_mem[377] = 16'b0000100001010000;
assign sigmoid_mem[378] = 16'b0000100001011100;
assign sigmoid_mem[379] = 16'b0000100001101001;
assign sigmoid_mem[380] = 16'b0000100001110101;
assign sigmoid_mem[381] = 16'b0000100010000010;
assign sigmoid_mem[382] = 16'b0000100010001110;
assign sigmoid_mem[383] = 16'b0000100010011011;
assign sigmoid_mem[384] = 16'b0000100010100111;
assign sigmoid_mem[385] = 16'b0000100010110100;
assign sigmoid_mem[386] = 16'b0000100011000001;
assign sigmoid_mem[387] = 16'b0000100011001101;
assign sigmoid_mem[388] = 16'b0000100011011010;
assign sigmoid_mem[389] = 16'b0000100011100111;
assign sigmoid_mem[390] = 16'b0000100011110100;
assign sigmoid_mem[391] = 16'b0000100100000001;
assign sigmoid_mem[392] = 16'b0000100100001110;
assign sigmoid_mem[393] = 16'b0000100100011011;
assign sigmoid_mem[394] = 16'b0000100100101000;
assign sigmoid_mem[395] = 16'b0000100100110101;
assign sigmoid_mem[396] = 16'b0000100101000010;
assign sigmoid_mem[397] = 16'b0000100101001111;
assign sigmoid_mem[398] = 16'b0000100101011100;
assign sigmoid_mem[399] = 16'b0000100101101010;
assign sigmoid_mem[400] = 16'b0000100101110111;
assign sigmoid_mem[401] = 16'b0000100110000100;
assign sigmoid_mem[402] = 16'b0000100110010010;
assign sigmoid_mem[403] = 16'b0000100110011111;
assign sigmoid_mem[404] = 16'b0000100110101101;
assign sigmoid_mem[405] = 16'b0000100110111010;
assign sigmoid_mem[406] = 16'b0000100111001000;
assign sigmoid_mem[407] = 16'b0000100111010101;
assign sigmoid_mem[408] = 16'b0000100111100011;
assign sigmoid_mem[409] = 16'b0000100111110001;
assign sigmoid_mem[410] = 16'b0000100111111110;
assign sigmoid_mem[411] = 16'b0000101000001100;
assign sigmoid_mem[412] = 16'b0000101000011010;
assign sigmoid_mem[413] = 16'b0000101000101000;
assign sigmoid_mem[414] = 16'b0000101000110110;
assign sigmoid_mem[415] = 16'b0000101001000100;
assign sigmoid_mem[416] = 16'b0000101001010010;
assign sigmoid_mem[417] = 16'b0000101001100000;
assign sigmoid_mem[418] = 16'b0000101001101110;
assign sigmoid_mem[419] = 16'b0000101001111100;
assign sigmoid_mem[420] = 16'b0000101010001010;
assign sigmoid_mem[421] = 16'b0000101010011000;
assign sigmoid_mem[422] = 16'b0000101010100110;
assign sigmoid_mem[423] = 16'b0000101010110100;
assign sigmoid_mem[424] = 16'b0000101011000011;
assign sigmoid_mem[425] = 16'b0000101011010001;
assign sigmoid_mem[426] = 16'b0000101011011111;
assign sigmoid_mem[427] = 16'b0000101011101110;
assign sigmoid_mem[428] = 16'b0000101011111100;
assign sigmoid_mem[429] = 16'b0000101100001011;
assign sigmoid_mem[430] = 16'b0000101100011001;
assign sigmoid_mem[431] = 16'b0000101100101000;
assign sigmoid_mem[432] = 16'b0000101100110110;
assign sigmoid_mem[433] = 16'b0000101101000101;
assign sigmoid_mem[434] = 16'b0000101101010011;
assign sigmoid_mem[435] = 16'b0000101101100010;
assign sigmoid_mem[436] = 16'b0000101101110001;
assign sigmoid_mem[437] = 16'b0000101101111111;
assign sigmoid_mem[438] = 16'b0000101110001110;
assign sigmoid_mem[439] = 16'b0000101110011101;
assign sigmoid_mem[440] = 16'b0000101110101100;
assign sigmoid_mem[441] = 16'b0000101110111011;
assign sigmoid_mem[442] = 16'b0000101111001001;
assign sigmoid_mem[443] = 16'b0000101111011000;
assign sigmoid_mem[444] = 16'b0000101111100111;
assign sigmoid_mem[445] = 16'b0000101111110110;
assign sigmoid_mem[446] = 16'b0000110000000101;
assign sigmoid_mem[447] = 16'b0000110000010100;
assign sigmoid_mem[448] = 16'b0000110000100011;
assign sigmoid_mem[449] = 16'b0000110000110010;
assign sigmoid_mem[450] = 16'b0000110001000010;
assign sigmoid_mem[451] = 16'b0000110001010001;
assign sigmoid_mem[452] = 16'b0000110001100000;
assign sigmoid_mem[453] = 16'b0000110001101111;
assign sigmoid_mem[454] = 16'b0000110001111110;
assign sigmoid_mem[455] = 16'b0000110010001110;
assign sigmoid_mem[456] = 16'b0000110010011101;
assign sigmoid_mem[457] = 16'b0000110010101100;
assign sigmoid_mem[458] = 16'b0000110010111011;
assign sigmoid_mem[459] = 16'b0000110011001011;
assign sigmoid_mem[460] = 16'b0000110011011010;
assign sigmoid_mem[461] = 16'b0000110011101010;
assign sigmoid_mem[462] = 16'b0000110011111001;
assign sigmoid_mem[463] = 16'b0000110100001000;
assign sigmoid_mem[464] = 16'b0000110100011000;
assign sigmoid_mem[465] = 16'b0000110100100111;
assign sigmoid_mem[466] = 16'b0000110100110111;
assign sigmoid_mem[467] = 16'b0000110101000110;
assign sigmoid_mem[468] = 16'b0000110101010110;
assign sigmoid_mem[469] = 16'b0000110101100101;
assign sigmoid_mem[470] = 16'b0000110101110101;
assign sigmoid_mem[471] = 16'b0000110110000101;
assign sigmoid_mem[472] = 16'b0000110110010100;
assign sigmoid_mem[473] = 16'b0000110110100100;
assign sigmoid_mem[474] = 16'b0000110110110100;
assign sigmoid_mem[475] = 16'b0000110111000011;
assign sigmoid_mem[476] = 16'b0000110111010011;
assign sigmoid_mem[477] = 16'b0000110111100011;
assign sigmoid_mem[478] = 16'b0000110111110010;
assign sigmoid_mem[479] = 16'b0000111000000010;
assign sigmoid_mem[480] = 16'b0000111000010010;
assign sigmoid_mem[481] = 16'b0000111000100010;
assign sigmoid_mem[482] = 16'b0000111000110001;
assign sigmoid_mem[483] = 16'b0000111001000001;
assign sigmoid_mem[484] = 16'b0000111001010001;
assign sigmoid_mem[485] = 16'b0000111001100001;
assign sigmoid_mem[486] = 16'b0000111001110001;
assign sigmoid_mem[487] = 16'b0000111010000001;
assign sigmoid_mem[488] = 16'b0000111010010000;
assign sigmoid_mem[489] = 16'b0000111010100000;
assign sigmoid_mem[490] = 16'b0000111010110000;
assign sigmoid_mem[491] = 16'b0000111011000000;
assign sigmoid_mem[492] = 16'b0000111011010000;
assign sigmoid_mem[493] = 16'b0000111011100000;
assign sigmoid_mem[494] = 16'b0000111011110000;
assign sigmoid_mem[495] = 16'b0000111100000000;
assign sigmoid_mem[496] = 16'b0000111100010000;
assign sigmoid_mem[497] = 16'b0000111100100000;
assign sigmoid_mem[498] = 16'b0000111100110000;
assign sigmoid_mem[499] = 16'b0000111101000000;
assign sigmoid_mem[500] = 16'b0000111101010000;
assign sigmoid_mem[501] = 16'b0000111101100000;
assign sigmoid_mem[502] = 16'b0000111101110000;
assign sigmoid_mem[503] = 16'b0000111110000000;
assign sigmoid_mem[504] = 16'b0000111110010000;
assign sigmoid_mem[505] = 16'b0000111110100000;
assign sigmoid_mem[506] = 16'b0000111110110000;
assign sigmoid_mem[507] = 16'b0000111111000000;
assign sigmoid_mem[508] = 16'b0000111111010000;
assign sigmoid_mem[509] = 16'b0000111111100000;
assign sigmoid_mem[510] = 16'b0000111111110000;
assign sigmoid_mem[511] = 16'b0001000000000000;
assign sigmoid_mem[512] = 16'b0001000000001111;
assign sigmoid_mem[513] = 16'b0001000000011111;
assign sigmoid_mem[514] = 16'b0001000000101111;
assign sigmoid_mem[515] = 16'b0001000000111111;
assign sigmoid_mem[516] = 16'b0001000001001111;
assign sigmoid_mem[517] = 16'b0001000001011111;
assign sigmoid_mem[518] = 16'b0001000001101111;
assign sigmoid_mem[519] = 16'b0001000001111111;
assign sigmoid_mem[520] = 16'b0001000010001111;
assign sigmoid_mem[521] = 16'b0001000010011111;
assign sigmoid_mem[522] = 16'b0001000010101111;
assign sigmoid_mem[523] = 16'b0001000010111111;
assign sigmoid_mem[524] = 16'b0001000011001111;
assign sigmoid_mem[525] = 16'b0001000011011111;
assign sigmoid_mem[526] = 16'b0001000011101111;
assign sigmoid_mem[527] = 16'b0001000011111111;
assign sigmoid_mem[528] = 16'b0001000100001111;
assign sigmoid_mem[529] = 16'b0001000100011111;
assign sigmoid_mem[530] = 16'b0001000100101111;
assign sigmoid_mem[531] = 16'b0001000100111111;
assign sigmoid_mem[532] = 16'b0001000101001111;
assign sigmoid_mem[533] = 16'b0001000101011111;
assign sigmoid_mem[534] = 16'b0001000101101111;
assign sigmoid_mem[535] = 16'b0001000101111110;
assign sigmoid_mem[536] = 16'b0001000110001110;
assign sigmoid_mem[537] = 16'b0001000110011110;
assign sigmoid_mem[538] = 16'b0001000110101110;
assign sigmoid_mem[539] = 16'b0001000110111110;
assign sigmoid_mem[540] = 16'b0001000111001110;
assign sigmoid_mem[541] = 16'b0001000111011101;
assign sigmoid_mem[542] = 16'b0001000111101101;
assign sigmoid_mem[543] = 16'b0001000111111101;
assign sigmoid_mem[544] = 16'b0001001000001101;
assign sigmoid_mem[545] = 16'b0001001000011100;
assign sigmoid_mem[546] = 16'b0001001000101100;
assign sigmoid_mem[547] = 16'b0001001000111100;
assign sigmoid_mem[548] = 16'b0001001001001011;
assign sigmoid_mem[549] = 16'b0001001001011011;
assign sigmoid_mem[550] = 16'b0001001001101011;
assign sigmoid_mem[551] = 16'b0001001001111010;
assign sigmoid_mem[552] = 16'b0001001010001010;
assign sigmoid_mem[553] = 16'b0001001010011010;
assign sigmoid_mem[554] = 16'b0001001010101001;
assign sigmoid_mem[555] = 16'b0001001010111001;
assign sigmoid_mem[556] = 16'b0001001011001000;
assign sigmoid_mem[557] = 16'b0001001011011000;
assign sigmoid_mem[558] = 16'b0001001011100111;
assign sigmoid_mem[559] = 16'b0001001011110111;
assign sigmoid_mem[560] = 16'b0001001100000110;
assign sigmoid_mem[561] = 16'b0001001100010101;
assign sigmoid_mem[562] = 16'b0001001100100101;
assign sigmoid_mem[563] = 16'b0001001100110100;
assign sigmoid_mem[564] = 16'b0001001101000100;
assign sigmoid_mem[565] = 16'b0001001101010011;
assign sigmoid_mem[566] = 16'b0001001101100010;
assign sigmoid_mem[567] = 16'b0001001101110001;
assign sigmoid_mem[568] = 16'b0001001110000001;
assign sigmoid_mem[569] = 16'b0001001110010000;
assign sigmoid_mem[570] = 16'b0001001110011111;
assign sigmoid_mem[571] = 16'b0001001110101110;
assign sigmoid_mem[572] = 16'b0001001110111101;
assign sigmoid_mem[573] = 16'b0001001111001101;
assign sigmoid_mem[574] = 16'b0001001111011100;
assign sigmoid_mem[575] = 16'b0001001111101011;
assign sigmoid_mem[576] = 16'b0001001111111010;
assign sigmoid_mem[577] = 16'b0001010000001001;
assign sigmoid_mem[578] = 16'b0001010000011000;
assign sigmoid_mem[579] = 16'b0001010000100111;
assign sigmoid_mem[580] = 16'b0001010000110110;
assign sigmoid_mem[581] = 16'b0001010001000100;
assign sigmoid_mem[582] = 16'b0001010001010011;
assign sigmoid_mem[583] = 16'b0001010001100010;
assign sigmoid_mem[584] = 16'b0001010001110001;
assign sigmoid_mem[585] = 16'b0001010010000000;
assign sigmoid_mem[586] = 16'b0001010010001110;
assign sigmoid_mem[587] = 16'b0001010010011101;
assign sigmoid_mem[588] = 16'b0001010010101100;
assign sigmoid_mem[589] = 16'b0001010010111010;
assign sigmoid_mem[590] = 16'b0001010011001001;
assign sigmoid_mem[591] = 16'b0001010011010111;
assign sigmoid_mem[592] = 16'b0001010011100110;
assign sigmoid_mem[593] = 16'b0001010011110100;
assign sigmoid_mem[594] = 16'b0001010100000011;
assign sigmoid_mem[595] = 16'b0001010100010001;
assign sigmoid_mem[596] = 16'b0001010100100000;
assign sigmoid_mem[597] = 16'b0001010100101110;
assign sigmoid_mem[598] = 16'b0001010100111100;
assign sigmoid_mem[599] = 16'b0001010101001011;
assign sigmoid_mem[600] = 16'b0001010101011001;
assign sigmoid_mem[601] = 16'b0001010101100111;
assign sigmoid_mem[602] = 16'b0001010101110101;
assign sigmoid_mem[603] = 16'b0001010110000011;
assign sigmoid_mem[604] = 16'b0001010110010001;
assign sigmoid_mem[605] = 16'b0001010110011111;
assign sigmoid_mem[606] = 16'b0001010110101101;
assign sigmoid_mem[607] = 16'b0001010110111011;
assign sigmoid_mem[608] = 16'b0001010111001001;
assign sigmoid_mem[609] = 16'b0001010111010111;
assign sigmoid_mem[610] = 16'b0001010111100101;
assign sigmoid_mem[611] = 16'b0001010111110011;
assign sigmoid_mem[612] = 16'b0001011000000001;
assign sigmoid_mem[613] = 16'b0001011000001110;
assign sigmoid_mem[614] = 16'b0001011000011100;
assign sigmoid_mem[615] = 16'b0001011000101010;
assign sigmoid_mem[616] = 16'b0001011000110111;
assign sigmoid_mem[617] = 16'b0001011001000101;
assign sigmoid_mem[618] = 16'b0001011001010010;
assign sigmoid_mem[619] = 16'b0001011001100000;
assign sigmoid_mem[620] = 16'b0001011001101101;
assign sigmoid_mem[621] = 16'b0001011001111011;
assign sigmoid_mem[622] = 16'b0001011010001000;
assign sigmoid_mem[623] = 16'b0001011010010101;
assign sigmoid_mem[624] = 16'b0001011010100011;
assign sigmoid_mem[625] = 16'b0001011010110000;
assign sigmoid_mem[626] = 16'b0001011010111101;
assign sigmoid_mem[627] = 16'b0001011011001010;
assign sigmoid_mem[628] = 16'b0001011011010111;
assign sigmoid_mem[629] = 16'b0001011011100100;
assign sigmoid_mem[630] = 16'b0001011011110001;
assign sigmoid_mem[631] = 16'b0001011011111110;
assign sigmoid_mem[632] = 16'b0001011100001011;
assign sigmoid_mem[633] = 16'b0001011100011000;
assign sigmoid_mem[634] = 16'b0001011100100101;
assign sigmoid_mem[635] = 16'b0001011100110010;
assign sigmoid_mem[636] = 16'b0001011100111110;
assign sigmoid_mem[637] = 16'b0001011101001011;
assign sigmoid_mem[638] = 16'b0001011101011000;
assign sigmoid_mem[639] = 16'b0001011101100100;
assign sigmoid_mem[640] = 16'b0001011101110001;
assign sigmoid_mem[641] = 16'b0001011101111101;
assign sigmoid_mem[642] = 16'b0001011110001010;
assign sigmoid_mem[643] = 16'b0001011110010110;
assign sigmoid_mem[644] = 16'b0001011110100011;
assign sigmoid_mem[645] = 16'b0001011110101111;
assign sigmoid_mem[646] = 16'b0001011110111011;
assign sigmoid_mem[647] = 16'b0001011111001000;
assign sigmoid_mem[648] = 16'b0001011111010100;
assign sigmoid_mem[649] = 16'b0001011111100000;
assign sigmoid_mem[650] = 16'b0001011111101100;
assign sigmoid_mem[651] = 16'b0001011111111000;
assign sigmoid_mem[652] = 16'b0001100000000100;
assign sigmoid_mem[653] = 16'b0001100000010000;
assign sigmoid_mem[654] = 16'b0001100000011100;
assign sigmoid_mem[655] = 16'b0001100000101000;
assign sigmoid_mem[656] = 16'b0001100000110100;
assign sigmoid_mem[657] = 16'b0001100000111111;
assign sigmoid_mem[658] = 16'b0001100001001011;
assign sigmoid_mem[659] = 16'b0001100001010111;
assign sigmoid_mem[660] = 16'b0001100001100010;
assign sigmoid_mem[661] = 16'b0001100001101110;
assign sigmoid_mem[662] = 16'b0001100001111001;
assign sigmoid_mem[663] = 16'b0001100010000101;
assign sigmoid_mem[664] = 16'b0001100010010000;
assign sigmoid_mem[665] = 16'b0001100010011100;
assign sigmoid_mem[666] = 16'b0001100010100111;
assign sigmoid_mem[667] = 16'b0001100010110010;
assign sigmoid_mem[668] = 16'b0001100010111110;
assign sigmoid_mem[669] = 16'b0001100011001001;
assign sigmoid_mem[670] = 16'b0001100011010100;
assign sigmoid_mem[671] = 16'b0001100011011111;
assign sigmoid_mem[672] = 16'b0001100011101010;
assign sigmoid_mem[673] = 16'b0001100011110101;
assign sigmoid_mem[674] = 16'b0001100100000000;
assign sigmoid_mem[675] = 16'b0001100100001011;
assign sigmoid_mem[676] = 16'b0001100100010110;
assign sigmoid_mem[677] = 16'b0001100100100001;
assign sigmoid_mem[678] = 16'b0001100100101100;
assign sigmoid_mem[679] = 16'b0001100100110110;
assign sigmoid_mem[680] = 16'b0001100101000001;
assign sigmoid_mem[681] = 16'b0001100101001100;
assign sigmoid_mem[682] = 16'b0001100101010110;
assign sigmoid_mem[683] = 16'b0001100101100001;
assign sigmoid_mem[684] = 16'b0001100101101011;
assign sigmoid_mem[685] = 16'b0001100101110110;
assign sigmoid_mem[686] = 16'b0001100110000000;
assign sigmoid_mem[687] = 16'b0001100110001010;
assign sigmoid_mem[688] = 16'b0001100110010101;
assign sigmoid_mem[689] = 16'b0001100110011111;
assign sigmoid_mem[690] = 16'b0001100110101001;
assign sigmoid_mem[691] = 16'b0001100110110011;
assign sigmoid_mem[692] = 16'b0001100110111101;
assign sigmoid_mem[693] = 16'b0001100111000111;
assign sigmoid_mem[694] = 16'b0001100111010001;
assign sigmoid_mem[695] = 16'b0001100111011011;
assign sigmoid_mem[696] = 16'b0001100111100101;
assign sigmoid_mem[697] = 16'b0001100111101111;
assign sigmoid_mem[698] = 16'b0001100111111001;
assign sigmoid_mem[699] = 16'b0001101000000011;
assign sigmoid_mem[700] = 16'b0001101000001100;
assign sigmoid_mem[701] = 16'b0001101000010110;
assign sigmoid_mem[702] = 16'b0001101000100000;
assign sigmoid_mem[703] = 16'b0001101000101001;
assign sigmoid_mem[704] = 16'b0001101000110011;
assign sigmoid_mem[705] = 16'b0001101000111100;
assign sigmoid_mem[706] = 16'b0001101001000101;
assign sigmoid_mem[707] = 16'b0001101001001111;
assign sigmoid_mem[708] = 16'b0001101001011000;
assign sigmoid_mem[709] = 16'b0001101001100001;
assign sigmoid_mem[710] = 16'b0001101001101011;
assign sigmoid_mem[711] = 16'b0001101001110100;
assign sigmoid_mem[712] = 16'b0001101001111101;
assign sigmoid_mem[713] = 16'b0001101010000110;
assign sigmoid_mem[714] = 16'b0001101010001111;
assign sigmoid_mem[715] = 16'b0001101010011000;
assign sigmoid_mem[716] = 16'b0001101010100001;
assign sigmoid_mem[717] = 16'b0001101010101010;
assign sigmoid_mem[718] = 16'b0001101010110011;
assign sigmoid_mem[719] = 16'b0001101010111100;
assign sigmoid_mem[720] = 16'b0001101011000101;
assign sigmoid_mem[721] = 16'b0001101011001101;
assign sigmoid_mem[722] = 16'b0001101011010110;
assign sigmoid_mem[723] = 16'b0001101011011111;
assign sigmoid_mem[724] = 16'b0001101011100111;
assign sigmoid_mem[725] = 16'b0001101011110000;
assign sigmoid_mem[726] = 16'b0001101011111000;
assign sigmoid_mem[727] = 16'b0001101100000001;
assign sigmoid_mem[728] = 16'b0001101100001001;
assign sigmoid_mem[729] = 16'b0001101100010001;
assign sigmoid_mem[730] = 16'b0001101100011010;
assign sigmoid_mem[731] = 16'b0001101100100010;
assign sigmoid_mem[732] = 16'b0001101100101010;
assign sigmoid_mem[733] = 16'b0001101100110010;
assign sigmoid_mem[734] = 16'b0001101100111011;
assign sigmoid_mem[735] = 16'b0001101101000011;
assign sigmoid_mem[736] = 16'b0001101101001011;
assign sigmoid_mem[737] = 16'b0001101101010011;
assign sigmoid_mem[738] = 16'b0001101101011011;
assign sigmoid_mem[739] = 16'b0001101101100011;
assign sigmoid_mem[740] = 16'b0001101101101011;
assign sigmoid_mem[741] = 16'b0001101101110010;
assign sigmoid_mem[742] = 16'b0001101101111010;
assign sigmoid_mem[743] = 16'b0001101110000010;
assign sigmoid_mem[744] = 16'b0001101110001010;
assign sigmoid_mem[745] = 16'b0001101110010001;
assign sigmoid_mem[746] = 16'b0001101110011001;
assign sigmoid_mem[747] = 16'b0001101110100000;
assign sigmoid_mem[748] = 16'b0001101110101000;
assign sigmoid_mem[749] = 16'b0001101110101111;
assign sigmoid_mem[750] = 16'b0001101110110111;
assign sigmoid_mem[751] = 16'b0001101110111110;
assign sigmoid_mem[752] = 16'b0001101111000110;
assign sigmoid_mem[753] = 16'b0001101111001101;
assign sigmoid_mem[754] = 16'b0001101111010100;
assign sigmoid_mem[755] = 16'b0001101111011011;
assign sigmoid_mem[756] = 16'b0001101111100011;
assign sigmoid_mem[757] = 16'b0001101111101010;
assign sigmoid_mem[758] = 16'b0001101111110001;
assign sigmoid_mem[759] = 16'b0001101111111000;
assign sigmoid_mem[760] = 16'b0001101111111111;
assign sigmoid_mem[761] = 16'b0001110000000110;
assign sigmoid_mem[762] = 16'b0001110000001101;
assign sigmoid_mem[763] = 16'b0001110000010100;
assign sigmoid_mem[764] = 16'b0001110000011011;
assign sigmoid_mem[765] = 16'b0001110000100001;
assign sigmoid_mem[766] = 16'b0001110000101000;
assign sigmoid_mem[767] = 16'b0001110000101111;
assign sigmoid_mem[768] = 16'b0001110000110110;
assign sigmoid_mem[769] = 16'b0001110000111100;
assign sigmoid_mem[770] = 16'b0001110001000011;
assign sigmoid_mem[771] = 16'b0001110001001010;
assign sigmoid_mem[772] = 16'b0001110001010000;
assign sigmoid_mem[773] = 16'b0001110001010111;
assign sigmoid_mem[774] = 16'b0001110001011101;
assign sigmoid_mem[775] = 16'b0001110001100011;
assign sigmoid_mem[776] = 16'b0001110001101010;
assign sigmoid_mem[777] = 16'b0001110001110000;
assign sigmoid_mem[778] = 16'b0001110001110111;
assign sigmoid_mem[779] = 16'b0001110001111101;
assign sigmoid_mem[780] = 16'b0001110010000011;
assign sigmoid_mem[781] = 16'b0001110010001001;
assign sigmoid_mem[782] = 16'b0001110010001111;
assign sigmoid_mem[783] = 16'b0001110010010101;
assign sigmoid_mem[784] = 16'b0001110010011100;
assign sigmoid_mem[785] = 16'b0001110010100010;
assign sigmoid_mem[786] = 16'b0001110010101000;
assign sigmoid_mem[787] = 16'b0001110010101110;
assign sigmoid_mem[788] = 16'b0001110010110100;
assign sigmoid_mem[789] = 16'b0001110010111001;
assign sigmoid_mem[790] = 16'b0001110010111111;
assign sigmoid_mem[791] = 16'b0001110011000101;
assign sigmoid_mem[792] = 16'b0001110011001011;
assign sigmoid_mem[793] = 16'b0001110011010001;
assign sigmoid_mem[794] = 16'b0001110011010110;
assign sigmoid_mem[795] = 16'b0001110011011100;
assign sigmoid_mem[796] = 16'b0001110011100010;
assign sigmoid_mem[797] = 16'b0001110011100111;
assign sigmoid_mem[798] = 16'b0001110011101101;
assign sigmoid_mem[799] = 16'b0001110011110010;
assign sigmoid_mem[800] = 16'b0001110011111000;
assign sigmoid_mem[801] = 16'b0001110011111101;
assign sigmoid_mem[802] = 16'b0001110100000011;
assign sigmoid_mem[803] = 16'b0001110100001000;
assign sigmoid_mem[804] = 16'b0001110100001110;
assign sigmoid_mem[805] = 16'b0001110100010011;
assign sigmoid_mem[806] = 16'b0001110100011000;
assign sigmoid_mem[807] = 16'b0001110100011101;
assign sigmoid_mem[808] = 16'b0001110100100011;
assign sigmoid_mem[809] = 16'b0001110100101000;
assign sigmoid_mem[810] = 16'b0001110100101101;
assign sigmoid_mem[811] = 16'b0001110100110010;
assign sigmoid_mem[812] = 16'b0001110100110111;
assign sigmoid_mem[813] = 16'b0001110100111100;
assign sigmoid_mem[814] = 16'b0001110101000001;
assign sigmoid_mem[815] = 16'b0001110101000110;
assign sigmoid_mem[816] = 16'b0001110101001011;
assign sigmoid_mem[817] = 16'b0001110101010000;
assign sigmoid_mem[818] = 16'b0001110101010101;
assign sigmoid_mem[819] = 16'b0001110101011010;
assign sigmoid_mem[820] = 16'b0001110101011111;
assign sigmoid_mem[821] = 16'b0001110101100100;
assign sigmoid_mem[822] = 16'b0001110101101000;
assign sigmoid_mem[823] = 16'b0001110101101101;
assign sigmoid_mem[824] = 16'b0001110101110010;
assign sigmoid_mem[825] = 16'b0001110101110111;
assign sigmoid_mem[826] = 16'b0001110101111011;
assign sigmoid_mem[827] = 16'b0001110110000000;
assign sigmoid_mem[828] = 16'b0001110110000100;
assign sigmoid_mem[829] = 16'b0001110110001001;
assign sigmoid_mem[830] = 16'b0001110110001110;
assign sigmoid_mem[831] = 16'b0001110110010010;
assign sigmoid_mem[832] = 16'b0001110110010111;
assign sigmoid_mem[833] = 16'b0001110110011011;
assign sigmoid_mem[834] = 16'b0001110110011111;
assign sigmoid_mem[835] = 16'b0001110110100100;
assign sigmoid_mem[836] = 16'b0001110110101000;
assign sigmoid_mem[837] = 16'b0001110110101100;
assign sigmoid_mem[838] = 16'b0001110110110001;
assign sigmoid_mem[839] = 16'b0001110110110101;
assign sigmoid_mem[840] = 16'b0001110110111001;
assign sigmoid_mem[841] = 16'b0001110110111101;
assign sigmoid_mem[842] = 16'b0001110111000010;
assign sigmoid_mem[843] = 16'b0001110111000110;
assign sigmoid_mem[844] = 16'b0001110111001010;
assign sigmoid_mem[845] = 16'b0001110111001110;
assign sigmoid_mem[846] = 16'b0001110111010010;
assign sigmoid_mem[847] = 16'b0001110111010110;
assign sigmoid_mem[848] = 16'b0001110111011010;
assign sigmoid_mem[849] = 16'b0001110111011110;
assign sigmoid_mem[850] = 16'b0001110111100010;
assign sigmoid_mem[851] = 16'b0001110111100110;
assign sigmoid_mem[852] = 16'b0001110111101010;
assign sigmoid_mem[853] = 16'b0001110111101110;
assign sigmoid_mem[854] = 16'b0001110111110010;
assign sigmoid_mem[855] = 16'b0001110111110110;
assign sigmoid_mem[856] = 16'b0001110111111001;
assign sigmoid_mem[857] = 16'b0001110111111101;
assign sigmoid_mem[858] = 16'b0001111000000001;
assign sigmoid_mem[859] = 16'b0001111000000101;
assign sigmoid_mem[860] = 16'b0001111000001000;
assign sigmoid_mem[861] = 16'b0001111000001100;
assign sigmoid_mem[862] = 16'b0001111000010000;
assign sigmoid_mem[863] = 16'b0001111000010011;
assign sigmoid_mem[864] = 16'b0001111000010111;
assign sigmoid_mem[865] = 16'b0001111000011010;
assign sigmoid_mem[866] = 16'b0001111000011110;
assign sigmoid_mem[867] = 16'b0001111000100010;
assign sigmoid_mem[868] = 16'b0001111000100101;
assign sigmoid_mem[869] = 16'b0001111000101001;
assign sigmoid_mem[870] = 16'b0001111000101100;
assign sigmoid_mem[871] = 16'b0001111000101111;
assign sigmoid_mem[872] = 16'b0001111000110011;
assign sigmoid_mem[873] = 16'b0001111000110110;
assign sigmoid_mem[874] = 16'b0001111000111010;
assign sigmoid_mem[875] = 16'b0001111000111101;
assign sigmoid_mem[876] = 16'b0001111001000000;
assign sigmoid_mem[877] = 16'b0001111001000100;
assign sigmoid_mem[878] = 16'b0001111001000111;
assign sigmoid_mem[879] = 16'b0001111001001010;
assign sigmoid_mem[880] = 16'b0001111001001101;
assign sigmoid_mem[881] = 16'b0001111001010000;
assign sigmoid_mem[882] = 16'b0001111001010100;
assign sigmoid_mem[883] = 16'b0001111001010111;
assign sigmoid_mem[884] = 16'b0001111001011010;
assign sigmoid_mem[885] = 16'b0001111001011101;
assign sigmoid_mem[886] = 16'b0001111001100000;
assign sigmoid_mem[887] = 16'b0001111001100011;
assign sigmoid_mem[888] = 16'b0001111001100110;
assign sigmoid_mem[889] = 16'b0001111001101001;
assign sigmoid_mem[890] = 16'b0001111001101100;
assign sigmoid_mem[891] = 16'b0001111001101111;
assign sigmoid_mem[892] = 16'b0001111001110010;
assign sigmoid_mem[893] = 16'b0001111001110101;
assign sigmoid_mem[894] = 16'b0001111001111000;
assign sigmoid_mem[895] = 16'b0001111001111011;
assign sigmoid_mem[896] = 16'b0001111001111110;
assign sigmoid_mem[897] = 16'b0001111010000001;
assign sigmoid_mem[898] = 16'b0001111010000100;
assign sigmoid_mem[899] = 16'b0001111010000110;
assign sigmoid_mem[900] = 16'b0001111010001001;
assign sigmoid_mem[901] = 16'b0001111010001100;
assign sigmoid_mem[902] = 16'b0001111010001111;
assign sigmoid_mem[903] = 16'b0001111010010001;
assign sigmoid_mem[904] = 16'b0001111010010100;
assign sigmoid_mem[905] = 16'b0001111010010111;
assign sigmoid_mem[906] = 16'b0001111010011010;
assign sigmoid_mem[907] = 16'b0001111010011100;
assign sigmoid_mem[908] = 16'b0001111010011111;
assign sigmoid_mem[909] = 16'b0001111010100010;
assign sigmoid_mem[910] = 16'b0001111010100100;
assign sigmoid_mem[911] = 16'b0001111010100111;
assign sigmoid_mem[912] = 16'b0001111010101001;
assign sigmoid_mem[913] = 16'b0001111010101100;
assign sigmoid_mem[914] = 16'b0001111010101110;
assign sigmoid_mem[915] = 16'b0001111010110001;
assign sigmoid_mem[916] = 16'b0001111010110011;
assign sigmoid_mem[917] = 16'b0001111010110110;
assign sigmoid_mem[918] = 16'b0001111010111000;
assign sigmoid_mem[919] = 16'b0001111010111011;
assign sigmoid_mem[920] = 16'b0001111010111101;
assign sigmoid_mem[921] = 16'b0001111011000000;
assign sigmoid_mem[922] = 16'b0001111011000010;
assign sigmoid_mem[923] = 16'b0001111011000100;
assign sigmoid_mem[924] = 16'b0001111011000111;
assign sigmoid_mem[925] = 16'b0001111011001001;
assign sigmoid_mem[926] = 16'b0001111011001011;
assign sigmoid_mem[927] = 16'b0001111011001110;
assign sigmoid_mem[928] = 16'b0001111011010000;
assign sigmoid_mem[929] = 16'b0001111011010010;
assign sigmoid_mem[930] = 16'b0001111011010101;
assign sigmoid_mem[931] = 16'b0001111011010111;
assign sigmoid_mem[932] = 16'b0001111011011001;
assign sigmoid_mem[933] = 16'b0001111011011011;
assign sigmoid_mem[934] = 16'b0001111011011101;
assign sigmoid_mem[935] = 16'b0001111011100000;
assign sigmoid_mem[936] = 16'b0001111011100010;
assign sigmoid_mem[937] = 16'b0001111011100100;
assign sigmoid_mem[938] = 16'b0001111011100110;
assign sigmoid_mem[939] = 16'b0001111011101000;
assign sigmoid_mem[940] = 16'b0001111011101010;
assign sigmoid_mem[941] = 16'b0001111011101100;
assign sigmoid_mem[942] = 16'b0001111011101110;
assign sigmoid_mem[943] = 16'b0001111011110000;
assign sigmoid_mem[944] = 16'b0001111011110010;
assign sigmoid_mem[945] = 16'b0001111011110101;
assign sigmoid_mem[946] = 16'b0001111011110111;
assign sigmoid_mem[947] = 16'b0001111011111001;
assign sigmoid_mem[948] = 16'b0001111011111011;
assign sigmoid_mem[949] = 16'b0001111011111100;
assign sigmoid_mem[950] = 16'b0001111011111110;
assign sigmoid_mem[951] = 16'b0001111100000000;
assign sigmoid_mem[952] = 16'b0001111100000010;
assign sigmoid_mem[953] = 16'b0001111100000100;
assign sigmoid_mem[954] = 16'b0001111100000110;
assign sigmoid_mem[955] = 16'b0001111100001000;
assign sigmoid_mem[956] = 16'b0001111100001010;
assign sigmoid_mem[957] = 16'b0001111100001100;
assign sigmoid_mem[958] = 16'b0001111100001110;
assign sigmoid_mem[959] = 16'b0001111100001111;
assign sigmoid_mem[960] = 16'b0001111100010001;
assign sigmoid_mem[961] = 16'b0001111100010011;
assign sigmoid_mem[962] = 16'b0001111100010101;
assign sigmoid_mem[963] = 16'b0001111100010111;
assign sigmoid_mem[964] = 16'b0001111100011000;
assign sigmoid_mem[965] = 16'b0001111100011010;
assign sigmoid_mem[966] = 16'b0001111100011100;
assign sigmoid_mem[967] = 16'b0001111100011110;
assign sigmoid_mem[968] = 16'b0001111100011111;
assign sigmoid_mem[969] = 16'b0001111100100001;
assign sigmoid_mem[970] = 16'b0001111100100011;
assign sigmoid_mem[971] = 16'b0001111100100100;
assign sigmoid_mem[972] = 16'b0001111100100110;
assign sigmoid_mem[973] = 16'b0001111100101000;
assign sigmoid_mem[974] = 16'b0001111100101001;
assign sigmoid_mem[975] = 16'b0001111100101011;
assign sigmoid_mem[976] = 16'b0001111100101100;
assign sigmoid_mem[977] = 16'b0001111100101110;
assign sigmoid_mem[978] = 16'b0001111100110000;
assign sigmoid_mem[979] = 16'b0001111100110001;
assign sigmoid_mem[980] = 16'b0001111100110011;
assign sigmoid_mem[981] = 16'b0001111100110100;
assign sigmoid_mem[982] = 16'b0001111100110110;
assign sigmoid_mem[983] = 16'b0001111100110111;
assign sigmoid_mem[984] = 16'b0001111100111001;
assign sigmoid_mem[985] = 16'b0001111100111010;
assign sigmoid_mem[986] = 16'b0001111100111100;
assign sigmoid_mem[987] = 16'b0001111100111101;
assign sigmoid_mem[988] = 16'b0001111100111111;
assign sigmoid_mem[989] = 16'b0001111101000000;
assign sigmoid_mem[990] = 16'b0001111101000010;
assign sigmoid_mem[991] = 16'b0001111101000011;
assign sigmoid_mem[992] = 16'b0001111101000101;
assign sigmoid_mem[993] = 16'b0001111101000110;
assign sigmoid_mem[994] = 16'b0001111101001000;
assign sigmoid_mem[995] = 16'b0001111101001001;
assign sigmoid_mem[996] = 16'b0001111101001010;
assign sigmoid_mem[997] = 16'b0001111101001100;
assign sigmoid_mem[998] = 16'b0001111101001101;
assign sigmoid_mem[999] = 16'b0001111101001110;
assign sigmoid_mem[1000] = 16'b0001111101010000;
assign sigmoid_mem[1001] = 16'b0001111101010001;
assign sigmoid_mem[1002] = 16'b0001111101010010;
assign sigmoid_mem[1003] = 16'b0001111101010100;
assign sigmoid_mem[1004] = 16'b0001111101010101;
assign sigmoid_mem[1005] = 16'b0001111101010110;
assign sigmoid_mem[1006] = 16'b0001111101011000;
assign sigmoid_mem[1007] = 16'b0001111101011001;
assign sigmoid_mem[1008] = 16'b0001111101011010;
assign sigmoid_mem[1009] = 16'b0001111101011011;
assign sigmoid_mem[1010] = 16'b0001111101011101;
assign sigmoid_mem[1011] = 16'b0001111101011110;
assign sigmoid_mem[1012] = 16'b0001111101011111;
assign sigmoid_mem[1013] = 16'b0001111101100000;
assign sigmoid_mem[1014] = 16'b0001111101100010;
assign sigmoid_mem[1015] = 16'b0001111101100011;
assign sigmoid_mem[1016] = 16'b0001111101100100;
assign sigmoid_mem[1017] = 16'b0001111101100101;
assign sigmoid_mem[1018] = 16'b0001111101100110;
assign sigmoid_mem[1019] = 16'b0001111101101000;
assign sigmoid_mem[1020] = 16'b0001111101101001;
assign sigmoid_mem[1021] = 16'b0001111101101010;
assign sigmoid_mem[1022] = 16'b0001111101101011;
assign sigmoid_mem[1023] = 16'b1;
// ---------- End of AUTOGENERATED CODE -------------------- //

always @(posedge clk)
begin
    if($signed(x_trunc) >= 0)
        y <= x_trunc+(2**(MEM_SIZE-1));
    else 
        y <= x_trunc-(2**(MEM_SIZE-1));      
end

assign sigmoid_out = sigmoid_mem[y];

endmodule